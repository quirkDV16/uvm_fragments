module tb_top;

 import uvm_pkg::*;

  initial begin
    run_test("my_test");
  end
endmodule
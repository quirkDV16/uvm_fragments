import uvm_pkg::*;

`include "uvm_macros.svh"
`include "my_agent.sv"
`include "my_env.sv"
`include "my_test.sv"


module top;

int top_int;

initial run_test();

endmodule

module top;

  import uvm_pkg::*;
  //import pkg::*;

  initial
    run_test("test");
  
endmodule


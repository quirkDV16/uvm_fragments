module top();
 import uvm_pkg::*;
  initial begin
    run_test();
  end
endmodule : top



module top();

import test_pkg::*;
import uvm_pkg::*;


`include "uvm_macros.svh"

initial run_test("my_test");

endmodule
